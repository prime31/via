module sdl2
import via.libs.sdl2.c

pub const ( version = c.version )
