module tilemap


