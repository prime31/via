module c


pub struct C.FMOD_STUDIO_SYSTEM {}
pub struct C.FMOD_STUDIO_EVENTDESCRIPTION {}
pub struct C.FMOD_STUDIO_EVENTINSTANCE {}
pub struct C.FMOD_STUDIO_BUS {}
pub struct C.FMOD_STUDIO_VCA {}
pub struct C.FMOD_STUDIO_BANK {}
pub struct C.FMOD_STUDIO_COMMANDREPLAY {}
pub struct C.FMOD_STUDIO_BANK_INFO {}
pub struct C.FMOD_STUDIO_PARAMETER_ID {}
pub struct C.FMOD_STUDIO_PARAMETER_DESCRIPTION {}
pub struct C.FMOD_STUDIO_USER_PROPERTY {}
pub struct C.FMOD_STUDIO_PROGRAMMER_SOUND_PROPERTIES {}
pub struct C.FMOD_STUDIO_PLUGIN_INSTANCE_PROPERTIES {}
pub struct C.FMOD_STUDIO_TIMELINE_MARKER_PROPERTIES {}
pub struct C.FMOD_STUDIO_TIMELINE_BEAT_PROPERTIES {}
pub struct C.FMOD_STUDIO_ADVANCEDSETTINGS {}
pub struct C.FMOD_STUDIO_CPU_USAGE {}
pub struct C.FMOD_STUDIO_BUFFER_INFO {}
pub struct C.FMOD_STUDIO_BUFFER_USAGE {}
pub struct C.FMOD_STUDIO_SOUND_INFO {}
pub struct C.FMOD_STUDIO_COMMAND_INFO {}

