module core

pub struct SoundGroup {
pub:
	group &FMOD_SOUNDGROUP
}