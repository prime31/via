module core

pub struct Dsp {
pub:
	dsp &C.FMOD_DSP
}