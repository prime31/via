module sokol
import via.libs.flextgl

const (
	used_import0 = flextgl.used_import
)