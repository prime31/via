module core

pub struct SoundGroup {
pub:
	group &C.FMOD_SOUNDGROUP
}