module sokol

// TODO: why is this needed all of a sudden for macos to compile?
#include <OpenGL/gl3.h>