module core

pub struct Dsp {
pub:
	dsp &FMOD_DSP
}