module c

pub const ( used_import = 1 )

pub struct C.FMOD_SYSTEM {}
pub struct C.FMOD_SOUND {}
pub struct C.FMOD_CHANNELCONTROL {}
pub struct C.FMOD_CHANNEL {}
pub struct C.FMOD_CHANNELGROUP {}
pub struct C.FMOD_SOUNDGROUP {}
pub struct C.FMOD_REVERB3D {}
pub struct C.FMOD_DSP {}
pub struct C.FMOD_DSPCONNECTION {}
pub struct C.FMOD_POLYGON {}
pub struct C.FMOD_GEOMETRY {}
pub struct C.FMOD_SYNCPOINT {}
pub struct C.FMOD_ASYNCREADINFO {}
pub struct C.FMOD_VECTOR {}
pub struct C.FMOD_3D_ATTRIBUTES {}
pub struct C.FMOD_GUID {}
pub struct C.FMOD_PLUGINLIST {}
pub struct C.FMOD_ADVANCEDSETTINGS {}
pub struct C.FMOD_TAG {}
pub struct C.FMOD_CREATESOUNDEXINFO {}
pub struct C.FMOD_REVERB_PROPERTIES {}
pub struct C.FMOD_ERRORCALLBACK_INFO {}

